class yapp_tx_sequencer extends uvm_sequencer #(yapp_packet);

//parameterization creates a yapp_packet object handle req automatically which can be used

//component utility macro
`uvm_component_utils(yapp_tx_sequencer)
 
 //component constructor
 function new(string name, uvm_component parent);
	super.new(name, parent);
 endfunction
 
endclass